`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:00:36 10/17/2016 
// Design Name: 
// Module Name:    core 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module core(
    input hit,
    input clr,
    output [3:0] NOM,
    output [1:0] BIT,
    output [3:0] LE,
    output TX
    );
wire [3:0] rg_a;
//wire ;



endmodule
